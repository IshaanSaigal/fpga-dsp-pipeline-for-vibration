`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.06.2025 17:47:01
// Design Name: 
// Module Name: fft_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fft_top (
    input wire CLK100MHZ,       // 100MHz clock pin, Pin W5
    input wire RESET_N,         // Active-low reset switch, Pin R2
    
    inout wire MPU_SCL,         // PMOD JA, Pin J1
    inout wire MPU_SDA,         // PMOD JA, Pin L2
    // NOTE: Since both SDA and SCL (clock stretching) can be controlled by both i2c_master and slave (MPU6050),
    // these must be modelled as inout ports.
    
    output wire UART_TXD        // UART Transmit Data line, Pin A18
);
    
    // --- Internal Signals ---
    logic rst_n;                        // Internal active-low reset signal
    assign rst_n = RESET_N;
    // The above code seems redundant for the i2c_master and uart_tx modules, which both have active-low resets.
    // However, in case any other module in the future requires a reset signal, which may be active-high, we need to have the
    // wire rst_n which we can alter as per our requirements (active-high vs active-low), while still using the same external switch.
    
    
    // --- Internal Signals for I2C ---
    logic i2c_enable_to_master_reg;
    logic i2c_read_write_to_master_reg;
    logic [7:0] i2c_mosi_data_to_master_reg;
    logic [7:0] i2c_register_address_to_master_reg;
    localparam IC_MPU_DEVICE_ADDRESS = 7'h68;       // MPU-6050's I2C address. Since this is constant, we use localparam
    localparam I2C_CLK_DIVIDER = 16'd249;           // For 100kHz Standard Mode I2C. 16-bit to match i2c_master. Since this is constant, we use localparam
    // For 100MHz system clk, 100kHz SCL clk:
    // f_SCL = f_CLK / (4 * (divider + 1))
    // => 100kHz = 100MHz / (4 * (divider + 1))
    // => divider = 249
    
    logic [7:0] i2c_miso_data_from_master;
    logic i2c_busy_from_master;
    
    
    // --- Internal Signals for I2C burst read ---
    // NOTE: Having separate signals for the burst instance is recommended to avoid contention.
    // For example, we don't want the same enable signal for both the instances, otherwise they both might try to seize the bus at the same time.
    logic i2c_enable_burst_to_master_reg;
    logic i2c_read_write_burst_to_master_reg;
    logic [15:0] i2c_mosi_data_burst_to_master_reg;     // Only needed for initialization; never actually used since we never do burst writes
    logic [7:0] i2c_register_address_burst_to_master_reg;
    // NOTE: The localparams remain same as the single-byte i2c_master instance
    
    logic [15:0] i2c_miso_data_burst_from_master;       // For 16-bit accelerometer readings
    logic i2c_busy_burst_from_master;
    
    
    // --- Internal Signals for UART ---
    logic uart_tx_en_pulse_sig;         // 1-cycle enable pulse for UART TX module
    logic [7:0] data_to_transmit_reg;   // Register to hold the data to be sent
    
    logic uart_busy_sig;                // Busy signal from UART TX module
    
    
    // --- Internal Signals for Input FIFO Buffer ---
    logic           fifo_sync_reset;     // wire
    logic           reset_sync_reg1;
    logic           reset_sync_reg2;
    // The "srst" port of the FIFO Generator IP is a synchronous reset.
    // "Synchronous" means that the reset only happens on the rising edge of the clk.
    // We cannot directly connect to RESETN switch since that is asynchronous, and could cause metastability in the FIFO core.
    // Thus, we update this in a separate always_ff block, synchronised with the clk.
    // For this, we will use a two-flop synchronizer chain:
    always_ff @(posedge CLK100MHZ) begin
        // First flop: Samples the asynchronous switch input.
        // This flop is allowed to go metastable.
        // We also invert the signal here since your switch is active-low (rst_n).
        reset_sync_reg1 <= !rst_n; 
        
        // Second flop: Samples the output of the first flop.
        // It has a full clock cycle for the first flop to settle.
        // The output of this flop is guaranteed to be stable.
        reset_sync_reg2 <= reset_sync_reg1;
    end
    assign fifo_sync_reset = reset_sync_reg2;
    
    logic           fifo_in_write_en_reg;
    logic [15:0]    fifo_in_write_data_reg;
    
    logic           fifo_in_read_en_reg;
    logic [15:0]    fifo_in_read_data;
    
    logic           fifo_in_full;
    logic           fifo_in_empty;
    
    // Counter for counting inputting exactly 1024 words in the FIFO buffer (1026 is the actual depth):
    logic [10:0]    fifo_in_write_counter_reg; // 11 bits, since I want to include 1024 as a comparison
    
    
    // --- Internal Signals for the FFT IP ---
    logic [31:0]    m_axis_data_tdata_reg;
    logic           m_axis_data_tvalid_reg;
    logic           m_axis_data_tready;
    logic           m_axis_data_tlast_reg;
    
    logic [31:0]    s_axis_data_tdata;
    logic           s_axis_data_tvalid;
    logic           s_axis_data_tready;
    logic           s_axis_data_tlast;
    
    logic [10:0]    flit_transfer_counter_reg;
    
    
    // --- Internal Signals for Output FIFO Buffer ---
    logic           fifo_out_write_en;
    //logic [31:0]    fifo_out_write_data_reg;  // using an extra reg here wastes a clock cycle; we can directly connect FFT IP's output
    
    logic           fifo_out_read_en_reg;
    logic [31:0]    fifo_out_read_data;
    
    logic           fifo_out_full;
    logic           fifo_out_empty;
    
    //NOTE: This buffer's input logic is combinational, but output is sequential. Might need to change the output??.
    // Combinational logic is needed for writing AXI4-Stream in a single clock cycle.
    
    // Counter for counting inputting exactly 1024 words in the FIFO buffer (1026 is the actual depth):
    //logic [10:0]    fifo_out_write_counter_reg; // 11 bits, since I want to include 1024 as a comparison
    // not needed because tlast signal
    
    
    // --- Instantiating I2C Master module ---
    i2c_master i2c_master_inst (
        .clock(CLK100MHZ),
        .reset_n(rst_n),
        .enable(i2c_enable_to_master_reg),
        .read_write(i2c_read_write_to_master_reg),
        .mosi_data(i2c_mosi_data_to_master_reg),
        .register_address(i2c_register_address_to_master_reg),
        .device_address(IC_MPU_DEVICE_ADDRESS),
        .divider(I2C_CLK_DIVIDER),
        
        .miso_data(i2c_miso_data_from_master),
        .busy(i2c_busy_from_master),
        
        .external_serial_data(MPU_SDA),
        .external_serial_clock(MPU_SCL)
    );
    
    
    // --- Instantiating I2C Master module for burst reads (for accelerometer readings) ---
    i2c_master #(
        .NUMBER_OF_DATA_BYTES(2)    // This parameter allows this instance to perform both burst reads and writes upto 2 bytes
    )
    i2c_master_burst_inst (
        .clock(CLK100MHZ),
        .reset_n(rst_n),
        .enable(i2c_enable_burst_to_master_reg),
        .read_write(i2c_read_write_burst_to_master_reg),
        .mosi_data(i2c_mosi_data_burst_to_master_reg),
        .register_address(i2c_register_address_burst_to_master_reg),
        .device_address(IC_MPU_DEVICE_ADDRESS),
        .divider(I2C_CLK_DIVIDER),
        
        .miso_data(i2c_miso_data_burst_from_master),
        .busy(i2c_busy_burst_from_master),
        
        .external_serial_data(MPU_SDA),
        .external_serial_clock(MPU_SCL)
    );
    
    
    // --- Instantiating UART TX Module ---
    uart_tx #(
        .BIT_RATE(115200),          // Baud rate
        .CLK_HZ(100_000_000),       // System clock frequency
        .PAYLOAD_BITS(8),           // Number of data bits
        .STOP_BITS(1)               // Number of stop bits
    ) uart_transmitter_inst (
        .clk(CLK100MHZ),                    // System clock
        .resetn(rst_n),                     // Active-low reset
        .uart_txd(UART_TXD),                // UART transmit data output pin
        .uart_tx_busy(uart_busy_sig),       // UART busy status output
        .uart_tx_en(uart_tx_en_pulse_sig),  // UART transmit enable (1-cycle pulse)
        .uart_tx_data(data_to_transmit_reg) // Data to be transmitted
    );
    
    
    // --- Instantiating Input FIFO Buffer IP ---
    fifo_buffer in_fifo_buffer_inst (
        .clk(CLK100MHZ),                // input wire clk
        .srst(fifo_sync_reset),      // input wire srst
        
        .din(fifo_in_write_data_reg),   // input wire [15 : 0] din
        .wr_en(fifo_in_write_en_reg),   // input wire wr_en
        
        .rd_en(fifo_in_read_en_reg),    // input wire rd_en
        .dout(fifo_in_read_data),       // output wire [15 : 0] dout
        
        .full(fifo_in_full),            // output wire full
        .empty(fifo_in_empty)           // output wire empty
    );
    
    
    // --- Instantiating the FFT IP ---
    fft_ip fft_ip_inst (
        .aclk(CLK100MHZ),                                                // input wire aclk
        .aclken(1'b1),                                            // input wire aclken
        .aresetn(rst_n),                                          // input wire aresetn
        
        // unconnected:
        .s_axis_config_tdata(16'b0),                  // input wire [15 : 0] s_axis_config_tdata
        .s_axis_config_tvalid(1'b0),                // input wire s_axis_config_tvalid
        .s_axis_config_tready(s_axis_config_tready),                // output wire s_axis_config_tready
        
        .s_axis_data_tdata(m_axis_data_tdata_reg),                      // input wire [31 : 0] s_axis_data_tdata
        .s_axis_data_tvalid(m_axis_data_tvalid_reg),                    // input wire s_axis_data_tvalid
        .s_axis_data_tready(m_axis_data_tready),                    // output wire s_axis_data_tready
        .s_axis_data_tlast(m_axis_data_tlast_reg),                      // input wire s_axis_data_tlast
        
        .m_axis_data_tdata(s_axis_data_tdata),                      // output wire [31 : 0] m_axis_data_tdata
        .m_axis_data_tvalid(s_axis_data_tvalid),                    // output wire m_axis_data_tvalid
        .m_axis_data_tready(s_axis_data_tready),                    // input wire m_axis_data_tready
        .m_axis_data_tlast(s_axis_data_tlast),                      // output wire m_axis_data_tlast
        
        // unconnected:
        .event_frame_started(event_frame_started),                  // output wire event_frame_started
        .event_tlast_unexpected(event_tlast_unexpected),            // output wire event_tlast_unexpected
        .event_tlast_missing(event_tlast_missing),                  // output wire event_tlast_missing
        .event_status_channel_halt(event_status_channel_halt),      // output wire event_status_channel_halt
        .event_data_in_channel_halt(event_data_in_channel_halt),    // output wire event_data_in_channel_halt
        .event_data_out_channel_halt(event_data_out_channel_halt)  // output wire event_data_out_channel_halt
    );
    
    
    // --- Instantiating Output FIFO Buffer IP ---
    fifo_generator_0 out_fifo_buffer_inst (
        .clk(CLK100MHZ),      // input wire clk
        .srst(fifo_sync_reset),    // input wire srst // using same signal as the input fifo buffer
        
        .din(s_axis_data_tdata),      // input wire [31 : 0] din
        .wr_en(fifo_out_write_en),  // input wire wr_en
        
        .rd_en(fifo_out_read_en_reg),  // input wire rd_en
        .dout(fifo_out_read_data),    // output wire [31 : 0] dout
        
        .full(fifo_out_full),    // output wire full
        .empty(fifo_out_empty)  // output wire empty
    );
    
    
    // --- Defining the FSM states ---
    typedef enum logic [5:0] {
        S_IDLE,
        
        // 1. Writing to PWR_MGMT_1 register
        S_I2C_PWR_MGMT_1_CONFIG,                    // Configure the inputs to the i2c_master module
        S_I2C_PWR_MGMT_1_WAIT_BEFORE_ENABLE,        // Ensure that the inputs are stable for 1 clock cycle
        S_I2C_PWR_MGMT_1_ENABLE,                    // Enable the i2c_master module
        S_I2C_PWR_MGMT_1_BUSY_HIGH_ENABLE_LOW,      // If busy is HIGH, pull enable LOW
        S_I2C_PWR_MGMT_1_WAIT_BUSY_LOW,             // Wait till i2c_master busy wire is LOW
        
        // 2. Writing to ACCEL_CONFIG register
        S_I2C_ACCEL_CONFIG_CONFIG,                  // Configure the inputs to the i2c_master module
        S_I2C_ACCEL_CONFIG_WAIT_BEFORE_ENABLE,      // Ensure that the inputs are stable for 1 clock cycle
        S_I2C_ACCEL_CONFIG_ENABLE,                  // Enable the i2c_master module
        S_I2C_ACCEL_CONFIG_BUSY_HIGH_ENABLE_LOW,    // If busy is HIGH, pull enable LOW
        S_I2C_ACCEL_CONFIG_WAIT_BUSY_LOW,           // Wait till i2c_master busy wire is LOW
        
        // 3. Reading ACCEL_XOUT_H and ACCEL_XOUT_L registers (burst read)
        S_I2C_ACCEL_XOUT_CONFIG,                    // Configure the inputs to the burst instance of the i2c_master module
        S_I2C_ACCEL_XOUT_WAIT_BEFORE_ENABLE,        // Ensure that the inputs are stable for 1 clock cycle
        S_I2C_ACCEL_XOUT_ENABLE,                    // Enable the burst instance of the i2c_master module
        S_I2C_ACCEL_XOUT_BUSY_HIGH_ENABLE_LOW,      // If busy is HIGH, pull enable LOW
        S_I2C_ACCEL_XOUT_WAIT_BUSY_LOW,             // Wait till i2c_master busy wire is LOW
        S_I2C_ACCEL_XOUT_READ_OUTPUT,               // Read the ACCEL_XOUT_H register (ACCEL_XOUT_L is still on the output wire of the burst instance)
                                                    // NEW: Read the ACCEL_XOUT_H and ACCEL_XOUT_L registers.
        
        // 4. Inputting accelerometer readings to FIFO buffer:
        S_FIFO_IN_WRITE_ENABLE,
        
        // 5. Sending ACCEL_XOUT_H over UART
        S_UART_ACCEL_XOUT_H_PULSE_ENABLE,       // Pulse the uart_tx enable wire for 1 system clock cycle
        S_UART_ACCEL_XOUT_H_WAIT_BUSY_LOW,      // Wait till the uart_tx busy wire is LOW
        
        // 6. Sending ACCEL_XOUT_L over UART
        S_UART_ACCEL_XOUT_L_LATCH,              // Latch the ACCEL_XOUT_L value to the uart_tx input data_to_transmit_reg (previously stored ACCEL_XOUT_H)
        S_UART_ACCEL_XOUT_L_PULSE_ENABLE,       // Pulse the uart_tx enable wire for 1 system clock cycle
        S_UART_ACCEL_XOUT_L_WAIT_BUSY_LOW,      // Wait till the uart_tx busy wire is LOW
        
        // 7. Reading WHO_AM_I register
        S_I2C_WHO_AM_I_CONFIG,                  // Configure the inputs to the i2c_master module
        S_I2C_WHO_AM_I_WAIT_BEFORE_ENABLE,      // Ensure that the inputs are stable for 1 clock cycle
        S_I2C_WHO_AM_I_ENABLE,                  // Enable the i2c_master module
        S_I2C_WHO_AM_I_BUSY_HIGH_ENABLE_LOW,    // If busy is HIGH, pull enable LOW
        S_I2C_WHO_AM_I_WAIT_BUSY_LOW,           // Wait till i2c_master busy wire is LOW
        S_I2C_WHO_AM_I_READ_OUTPUT,             // Read the WHO_AM_I register's value
        
        // 8. Sending WHO_AM_I over UART
        S_UART_WHO_AM_I_PULSE_ENABLE,           // Pulse the uart_tx enable wire for 1 system clock cycle
        S_UART_WHO_AM_I_WAIT_BUSY_LOW,          // Wait till the uart_tx busy wire is LOW
        
        // 9. Inputting the FIFO buffer's values to the FFT IP once we have collected 1024 samples:
        S_FFT_IN_CONFIG,
        S_FFT_IN_ASSERT_TVALID,
        
        // 10. Inputting FFT IP's output to FIFO buffer:
        //S_FFT_WAIT_TVALID, // wait till the output tvalid is high
        //S_FIFO_OUT_WRITE_CONFIG, // put the write data on the fifo din bus
        //S_FIFO_OUT_WRITE_ENABLE,
        S_FFT_WAIT_TLAST,
        
        // 11. Sending FIFO buffer's data over UART (real higher byte):
        S_UART_FIFO_OUT_H_LATCH,             // Latch the ACCEL_XOUT_H value to the uart_tx input data_to_transmit_reg
        S_UART_FIFO_OUT_H_PULSE_ENABLE,       // Pulse the uart_tx enable wire for 1 system clock cycle
        S_UART_FIFO_OUT_H_WAIT_BUSY_LOW,      // Wait till the uart_tx busy wire is LOW
        
        // 12. Sending FIFO buffer's data over UART (real lower byte):
        S_UART_FIFO_OUT_L_LATCH,              // Latch the ACCEL_XOUT_L value to the uart_tx input data_to_transmit_reg (previously stored ACCEL_XOUT_H)
        S_UART_FIFO_OUT_L_PULSE_ENABLE,       // Pulse the uart_tx enable wire for 1 system clock cycle
        S_UART_FIFO_OUT_L_WAIT_BUSY_LOW,      // Wait till the uart_tx busy wire is LOW
        
        S_DONE
    } main_state_t;
    
    main_state_t current_state, next_state;
    
    // NOTE: We need a separate always_ff block to update current_state. Otherwise, if we used the same always_ff block as the
    // rest of the sequential logic, the case(current_state) won't know which current_state to use: the one that just updated
    // vs one that was used in the previous cycle. This causes a Synthesis Error.
    always_ff @(posedge CLK100MHZ or negedge rst_n) begin
        if (!rst_n) begin
            current_state <= S_IDLE;
        end else begin
            current_state <= next_state;
        end
    end
    
    
    // --- FSM Sequential Logic ---
    // NOTE: The I2C logic is both sequential and combinational
    always_ff @(posedge CLK100MHZ or negedge rst_n) begin
        if (!rst_n) begin
            // Reset values for all registers controlled by this FSM
            i2c_enable_to_master_reg <= 1'b0;
            i2c_read_write_to_master_reg <= 1'b0;
            i2c_mosi_data_to_master_reg <= 8'h00;
            i2c_register_address_to_master_reg <= 8'h00;
            
            i2c_enable_burst_to_master_reg <= 1'b0;
            i2c_read_write_burst_to_master_reg <= 1'b0;
            i2c_mosi_data_burst_to_master_reg <= 16'b0;     // Always remains 0, since we never need to burst write
            i2c_register_address_burst_to_master_reg <= 8'h00;
            
            data_to_transmit_reg <= 8'h00;
            
            fifo_in_write_en_reg <= 1'b0;
            fifo_in_write_data_reg <= 16'b0;
            fifo_in_read_en_reg <= 1'b0;
            fifo_in_write_counter_reg <= 11'b0;
            
            m_axis_data_tdata_reg <= 32'b0;
            m_axis_data_tvalid_reg <= 1'b0;
            m_axis_data_tlast_reg <= 1'b0;
            //s_axis_data_tready_reg <= 1'b0;
            flit_transfer_counter_reg <= 11'b0;
            
            //fifo_out_write_en_reg <= 1'b0;
            //fifo_out_write_data_reg <= 32'b0;
            fifo_out_read_en_reg <= 1'b0;
            
        end else begin
            // Defaults:
            i2c_enable_to_master_reg <= 1'b0;
            i2c_enable_burst_to_master_reg <= 1'b0;
            // The rest of the I2C registers are held undefined/latched right now
            
            fifo_in_write_en_reg <= 1'b0;
            fifo_in_read_en_reg <= 1'b0;
            // The rest of the input FIFO IP registers are held undefined/latched right now.
            
            m_axis_data_tvalid_reg <= 1'b0;
            m_axis_data_tlast_reg <= 1'b0;
            //s_axis_data_tready_reg <= 1'b0;
            // The rest of the FFT IP registers are held undefined/latched right now.
            
            //fifo_out_write_en_reg <= 1'b0;
            fifo_out_read_en_reg <= 1'b0;
            // The rest of the output FIFO IP registers are held undefined/latched right now.
            
            case (current_state)
                
                // 1. Writing to PWR_MGMT_1 register
                
                S_I2C_PWR_MGMT_1_CONFIG: begin
                    i2c_read_write_to_master_reg <= 1'b0;           // For writing
                    i2c_mosi_data_to_master_reg <= 8'h01;           // 1) Wake up; 2) Gyro-referenced PLL as clock; 3). Leave temperature sensing enabled 
                    i2c_register_address_to_master_reg <= 8'h6B;    // Address of the PWR_MGMT_1 register
                end
                
                S_I2C_PWR_MGMT_1_ENABLE: begin
                    i2c_enable_to_master_reg <= 1'b1;
                end
                
                S_I2C_PWR_MGMT_1_BUSY_HIGH_ENABLE_LOW: begin
                    if (!i2c_busy_from_master)
                        i2c_enable_to_master_reg <= 1'b1;   // Keep enable high if busy is low
                    else
                        i2c_enable_to_master_reg <= 1'b0;   // Keep enable low if busy is high
                end
                
                
                // 2. Writing to ACCEL_CONFIG register
                
                S_I2C_ACCEL_CONFIG_CONFIG: begin
                    i2c_read_write_to_master_reg <= 1'b0;           // For writing
                    i2c_mosi_data_to_master_reg <= 8'h10;           // For configuring full-scale range of accelerometer as +-8g
                    i2c_register_address_to_master_reg <= 8'h1C;    // Address of the ACCEL_CONFIG register
                end
                
                S_I2C_ACCEL_CONFIG_ENABLE: begin
                    i2c_enable_to_master_reg <= 1'b1;
                end
                
                S_I2C_ACCEL_CONFIG_BUSY_HIGH_ENABLE_LOW: begin
                    if (!i2c_busy_from_master)
                        i2c_enable_to_master_reg <= 1'b1;   // Keep enable high if busy is low
                    else
                        i2c_enable_to_master_reg <= 1'b0;   // Keep enable low if busy is high
                end
                
                
                // 3. Reading ACCEL_XOUT_H and ACCEL_XOUT_L (burst read)
                
                S_I2C_ACCEL_XOUT_CONFIG: begin
                    i2c_read_write_burst_to_master_reg <= 1'b1;         // For reading (burst read 2 bytes)
                    i2c_mosi_data_burst_to_master_reg <= 16'h00;        // We want to read, not write. But we should still define this with a fixed value
                    i2c_register_address_burst_to_master_reg <= 8'h3B;  // Address of the ACCEL_XOUT_H register. Both this and ACCEL_XOUT_L are burst read
                end
                
                S_I2C_ACCEL_XOUT_ENABLE: begin
                    i2c_enable_burst_to_master_reg <= 1'b1;
                end
                
                S_I2C_ACCEL_XOUT_BUSY_HIGH_ENABLE_LOW: begin
                    if (!i2c_busy_burst_from_master)
                        i2c_enable_burst_to_master_reg <= 1'b1;     // Keep enable high if busy is low
                    else
                        i2c_enable_burst_to_master_reg <= 1'b0;     // Keep enable low if busy is high
                end
                
                S_I2C_ACCEL_XOUT_READ_OUTPUT: begin
                    // Actually read the i2c_master master
                    fifo_in_write_data_reg <= i2c_miso_data_burst_from_master;
                    
                    // For UART:
                    data_to_transmit_reg <= i2c_miso_data_burst_from_master[15:8];
                    // We read the ACCEL_XOUT_H byte right now.
                    // The ACCEL_XOUT_L still remains on the i2c_miso_data_burst_from_master line, which we read later.
                end
                
                
                // 4. Inputting accelerometer readings to FIFO buffer:
                
                S_FIFO_IN_WRITE_ENABLE: begin
                    if (!fifo_in_full) begin
                        // Write to the FIFO buffer only if it has less than 1024 words (and it is NOT full, which it won't be since actual depth is 1026):
                        fifo_in_write_en_reg <= 1'b1;
                    end
                    
                    // Increment the counter:
                    fifo_in_write_counter_reg <= fifo_in_write_counter_reg + 1;
                end
                
                
                // 6. Sending ACCEL_XOUT_L over UART
                
                S_UART_ACCEL_XOUT_L_LATCH: begin
                    // Latch the ACCEL_XOUT_L to uart_tx's data_to_transmit_reg (previously ACCEL_XOUT_H) for transmission
                    data_to_transmit_reg <= i2c_miso_data_burst_from_master[7:0];
                end
                
                
                // 7. Reading WHO_AM_I register
                
                S_I2C_WHO_AM_I_CONFIG: begin
                    i2c_read_write_to_master_reg <= 1'b1;           // For reading
                    i2c_mosi_data_to_master_reg <= 8'h00;           // We want to read, not write. But we should still define this with a fixed value
                    i2c_register_address_to_master_reg <= 8'h75;    // Address of the WHO_AM_I register
                end
                
                S_I2C_WHO_AM_I_ENABLE: begin
                    i2c_enable_to_master_reg <= 1'b1;
                end
                
                S_I2C_WHO_AM_I_BUSY_HIGH_ENABLE_LOW: begin
                    if (!i2c_busy_from_master)
                        i2c_enable_to_master_reg <= 1'b1;   // Keep enable high if busy is low
                    else
                        i2c_enable_to_master_reg <= 1'b0;   // Keep enable low if busy is high
                end
                
                S_I2C_WHO_AM_I_READ_OUTPUT: begin
                    // Actually read the i2c_master master
                    data_to_transmit_reg <= i2c_miso_data_from_master;      // 8'h68 (ASCII 'h') is the ideal return from WHO_AM_I
                end
                
                
                // 9.
                
                S_FFT_IN_CONFIG: begin
                    fifo_in_write_counter_reg <= 11'b0; //reset this counter
                    
                    if (!fifo_in_empty)
                        m_axis_data_tdata_reg <= {16'b0, fifo_in_read_data}; // concatenation
                    
                    // need to assert tlast depending on a counter here
                    if (flit_transfer_counter_reg == 1023) // // 1023 means 1023 flits have been transferred; 1024th (last) is left
                        m_axis_data_tlast_reg <= 1'b1;
                end
                
                S_FFT_IN_ASSERT_TVALID: begin
                    m_axis_data_tvalid_reg <= 1'b1;
                    
                    if (m_axis_data_tready && !fifo_in_empty) begin // means current word will be inputted to the FFT IP; we should go to the next word
                        // Assert read enable to request the next word
                        fifo_in_read_en_reg <= 1'b1; // read; output is available on the same clock cycle
                        
                        // increment counter indicating a flit transfer:
                        flit_transfer_counter_reg <= flit_transfer_counter_reg + 1;
                    end
                end
                
                
                // 10.
                
                /*S_FIFO_OUT_WRITE_CONFIG: begin
                    if (s_axis_data_tvalid)
                        fifo_out_write_data_reg <= s_axis_data_tdata;
                end
                
                S_FFT_WAIT_TLAST: begin
                    if (s_axis_data_tvalid && !fifo_out_full) begin
                        fifo_out_write_en_reg <= 1'b1;
                        
                        // tready:
                        s_axis_data_tready_reg <= 1'b1;     // tvalid is high; we are making tready high => flit transfer occurs on NEXT cycle
                    end
                end*/
                
                S_FFT_WAIT_TLAST: begin
                    flit_transfer_counter_reg <= 10'b0; //reset this counter
                end
                
                
                // 11. Sending FIFO buffer's data over UART (higher byte):
                
                S_UART_FIFO_OUT_H_LATCH: begin
                    if (!fifo_out_empty) begin
                        // Latch the higher byte to uart_tx's data_to_transmit_reg for transmission
                        data_to_transmit_reg <= fifo_out_read_data[15:8];
                    end
                end
                
                
                // 12. Sending FIFO buffer's data over UART (lower byte):
                S_UART_FIFO_OUT_L_LATCH: begin
                    if (!fifo_out_empty) begin
                        // Latch the lower byte to uart_tx's data_to_transmit_reg for transmission
                        data_to_transmit_reg <= fifo_out_read_data[7:0];
                        
                        // Assert read enable to request the next word
                        fifo_out_read_en_reg <= 1'b1; // read; output is available on the same clock cycle
                    end
                end
                
            endcase
        end
    end
    
    
    // --- FSM Combinational Logic ---
    // NOTE: The UART logic is fully combinational
    always_comb begin
        // Defaults:
        uart_tx_en_pulse_sig = 1'b0;    // When in any other state except S_UART_PULSE_ENABLE, uart_tx_en_pulse_sig is LOW by default
        
        next_state = current_state;     // By default, stay in current_state, unless explicitly mentioned in a case
        
        s_axis_data_tready = 1'b0;
        fifo_out_write_en = 1'b0;
        
        case (current_state)
            S_IDLE: begin
                next_state = S_I2C_PWR_MGMT_1_CONFIG;
            end
            
            
            // 1. Writing to PWR_MGMT_1 register
            
            S_I2C_PWR_MGMT_1_CONFIG: begin
                next_state = S_I2C_PWR_MGMT_1_WAIT_BEFORE_ENABLE;
            end
            
            S_I2C_PWR_MGMT_1_WAIT_BEFORE_ENABLE: begin
                // Wait 1 clock cycle for the configuration values to stabilize
                if (!i2c_busy_from_master) begin
                    next_state = S_I2C_PWR_MGMT_1_ENABLE;               // If I2C core is idle, proceed to enable it
                end else begin
                    next_state = S_I2C_PWR_MGMT_1_WAIT_BEFORE_ENABLE;   // Else, keep waiting
                end
            end
            
            S_I2C_PWR_MGMT_1_ENABLE: begin
                next_state = S_I2C_PWR_MGMT_1_BUSY_HIGH_ENABLE_LOW;
            end
            
            S_I2C_PWR_MGMT_1_BUSY_HIGH_ENABLE_LOW: begin
                // Wait till busy signal is HIGH to set enable signal LOW
                if (!i2c_enable_to_master_reg && i2c_busy_from_master)
                    next_state = S_I2C_PWR_MGMT_1_WAIT_BUSY_LOW;
                else
                    next_state = S_I2C_PWR_MGMT_1_BUSY_HIGH_ENABLE_LOW;
            end
            
            S_I2C_PWR_MGMT_1_WAIT_BUSY_LOW: begin
                // Wait till busy is LOW, which means I2C transaction is complete
                if (!i2c_busy_from_master)
                    next_state = S_I2C_ACCEL_CONFIG_CONFIG;
                else
                    next_state = S_I2C_PWR_MGMT_1_WAIT_BUSY_LOW;
            end
            
            
            // 2. Writing to ACCEL_CONFIG register
            
            S_I2C_ACCEL_CONFIG_CONFIG: begin
                next_state = S_I2C_ACCEL_CONFIG_WAIT_BEFORE_ENABLE;
            end
            
            S_I2C_ACCEL_CONFIG_WAIT_BEFORE_ENABLE: begin
                // Wait 1 clock cycle for the configuration values to stabilize
                if (!i2c_busy_from_master) begin
                    next_state = S_I2C_ACCEL_CONFIG_ENABLE;             // If I2C core is idle, proceed to enable it
                end else begin
                    next_state = S_I2C_ACCEL_CONFIG_WAIT_BEFORE_ENABLE; // Else, keep waiting
                end
            end
            
            S_I2C_ACCEL_CONFIG_ENABLE: begin
                next_state = S_I2C_ACCEL_CONFIG_BUSY_HIGH_ENABLE_LOW;
            end
            
            S_I2C_ACCEL_CONFIG_BUSY_HIGH_ENABLE_LOW: begin
                // Wait till busy signal is HIGH to set enable signal LOW
                if (!i2c_enable_to_master_reg && i2c_busy_from_master)
                    next_state = S_I2C_ACCEL_CONFIG_WAIT_BUSY_LOW;
                else
                    next_state = S_I2C_ACCEL_CONFIG_BUSY_HIGH_ENABLE_LOW;
            end
            
            S_I2C_ACCEL_CONFIG_WAIT_BUSY_LOW: begin
                // Wait till busy is LOW, which means I2C transaction is complete
                if (!i2c_busy_from_master)
                    next_state = S_I2C_ACCEL_XOUT_CONFIG;
                else
                    next_state = S_I2C_ACCEL_CONFIG_WAIT_BUSY_LOW;
            end
            
            
            // 3. Reading ACCEL_XOUT_H and ACCEL_XOUT_L (burst read)
            
            S_I2C_ACCEL_XOUT_CONFIG: begin
                next_state = S_I2C_ACCEL_XOUT_WAIT_BEFORE_ENABLE;
            end
            
            S_I2C_ACCEL_XOUT_WAIT_BEFORE_ENABLE: begin
                // Wait 1 clock cycle for the configuration values to stabilize
                if (!i2c_busy_burst_from_master) begin
                    next_state = S_I2C_ACCEL_XOUT_ENABLE;               // If I2C burst instance is idle, proceed to enable it
                end else begin
                    next_state = S_I2C_ACCEL_XOUT_WAIT_BEFORE_ENABLE;   // Else, keep waiting
                end
            end
            
            S_I2C_ACCEL_XOUT_ENABLE: begin
                next_state = S_I2C_ACCEL_XOUT_BUSY_HIGH_ENABLE_LOW;
            end
            
            S_I2C_ACCEL_XOUT_BUSY_HIGH_ENABLE_LOW: begin
                // Wait till busy signal is HIGH to set enable signal LOW
                if (!i2c_enable_burst_to_master_reg && i2c_busy_burst_from_master)
                    next_state = S_I2C_ACCEL_XOUT_WAIT_BUSY_LOW;
                else
                    next_state = S_I2C_ACCEL_XOUT_BUSY_HIGH_ENABLE_LOW;
            end
            
            S_I2C_ACCEL_XOUT_WAIT_BUSY_LOW: begin
                // Wait till busy is LOW, which means I2C transaction is complete
                if (!i2c_busy_burst_from_master)
                    next_state = S_I2C_ACCEL_XOUT_READ_OUTPUT;
                else
                    next_state = S_I2C_ACCEL_XOUT_WAIT_BUSY_LOW;
            end
            
            S_I2C_ACCEL_XOUT_READ_OUTPUT: begin
                next_state = S_FIFO_IN_WRITE_ENABLE;
            end
            
            
            // 4. Inputting accelerometer readings to FIFO buffer:
            
            S_FIFO_IN_WRITE_ENABLE: begin
                next_state = S_UART_ACCEL_XOUT_H_PULSE_ENABLE;
            end
            
            
            // 5. Sending ACCEL_XOUT_H over UART
            
            S_UART_ACCEL_XOUT_H_PULSE_ENABLE: begin
                uart_tx_en_pulse_sig = !uart_busy_sig && rst_n;         // HIGH only when the UART TX module is NOT busy and NOT in reset
                // uart_tx_en_pulse_sig is HIGH for 1 cycle, since the FSM states last 1 clock cycle each
                
                if (uart_tx_en_pulse_sig)
                    next_state = S_UART_ACCEL_XOUT_H_WAIT_BUSY_LOW;     // Only transition to the next state once enable signal is HIGH
                else
                    next_state = S_UART_ACCEL_XOUT_H_PULSE_ENABLE;
            end
            
            S_UART_ACCEL_XOUT_H_WAIT_BUSY_LOW: begin
                // Transition when UART TX module is not busy, else wait here till communication is finished
                if (!uart_busy_sig)
                    next_state = S_UART_ACCEL_XOUT_L_LATCH;
                else
                    next_state = S_UART_ACCEL_XOUT_H_WAIT_BUSY_LOW;
            end
            
            
            // 6. Sending ACCEL_XOUT_L over UART
            
            S_UART_ACCEL_XOUT_L_LATCH: begin
                // Just wait 1 clock cycle to latch the ACCEL_XOUT_L to uart_tx's data_to_transmit_reg
                next_state = S_UART_ACCEL_XOUT_L_PULSE_ENABLE;
            end
            
            S_UART_ACCEL_XOUT_L_PULSE_ENABLE: begin
                uart_tx_en_pulse_sig = !uart_busy_sig && rst_n;         // HIGH only when the UART TX module is NOT busy and NOT in reset
                // uart_tx_en_pulse_sig is HIGH for 1 cycle, since the FSM states last 1 clock cycle each
                
                if (uart_tx_en_pulse_sig)
                    next_state = S_UART_ACCEL_XOUT_L_WAIT_BUSY_LOW;     // Only transition to the next state once enable signal is HIGH
                else
                    next_state = S_UART_ACCEL_XOUT_L_PULSE_ENABLE;
            end
            
            S_UART_ACCEL_XOUT_L_WAIT_BUSY_LOW: begin
                // Transition when UART TX module is not busy, else wait here till communication is finished
                if (!uart_busy_sig)
                    next_state = S_I2C_WHO_AM_I_CONFIG;
                else
                    next_state = S_UART_ACCEL_XOUT_L_WAIT_BUSY_LOW;
            end
            
            
            // 7. Reading WHO_AM_I register
            
            S_I2C_WHO_AM_I_CONFIG: begin
                next_state = S_I2C_WHO_AM_I_WAIT_BEFORE_ENABLE;
            end
            
            S_I2C_WHO_AM_I_WAIT_BEFORE_ENABLE: begin
                // Wait 1 clock cycle for the configuration values to stabilize
                if (!i2c_busy_from_master) begin
                    next_state = S_I2C_WHO_AM_I_ENABLE;             // If I2C core is idle, proceed to enable it
                end else begin
                    next_state = S_I2C_WHO_AM_I_WAIT_BEFORE_ENABLE; // Else, keep waiting
                end
            end
            
            S_I2C_WHO_AM_I_ENABLE: begin
                next_state = S_I2C_WHO_AM_I_BUSY_HIGH_ENABLE_LOW;
            end
            
            S_I2C_WHO_AM_I_BUSY_HIGH_ENABLE_LOW: begin
                // Wait till busy signal is HIGH to set enable signal LOW
                if (!i2c_enable_to_master_reg && i2c_busy_from_master)
                    next_state = S_I2C_WHO_AM_I_WAIT_BUSY_LOW;
                else
                    next_state = S_I2C_WHO_AM_I_BUSY_HIGH_ENABLE_LOW;
            end
            
            S_I2C_WHO_AM_I_WAIT_BUSY_LOW: begin
                // Wait till busy is LOW, which means I2C transaction is complete
                if (!i2c_busy_from_master)
                    next_state = S_I2C_WHO_AM_I_READ_OUTPUT;
                else
                    next_state = S_I2C_WHO_AM_I_WAIT_BUSY_LOW;
            end
            
            S_I2C_WHO_AM_I_READ_OUTPUT: begin
                next_state = S_UART_WHO_AM_I_PULSE_ENABLE;
            end
            
            
            // 8. Sending WHO_AM_I over UART
            
            S_UART_WHO_AM_I_PULSE_ENABLE: begin
                uart_tx_en_pulse_sig = !uart_busy_sig && rst_n;     // HIGH only when the UART TX module is NOT busy and NOT in reset
                // uart_tx_en_pulse_sig is HIGH for 1 cycle, since the FSM states last 1 clock cycle each
                
                if (uart_tx_en_pulse_sig)
                    next_state = S_UART_WHO_AM_I_WAIT_BUSY_LOW;     // Only transition to the next state once enable signal is HIGH
                else
                    next_state = S_UART_WHO_AM_I_PULSE_ENABLE;
            end
            
            S_UART_WHO_AM_I_WAIT_BUSY_LOW: begin
                // Transition when UART TX module is not busy, else wait here till communication is finished
                if (!uart_busy_sig) begin
                    if (fifo_in_write_counter_reg == 1024 || fifo_in_full) // go to fifo reading if counter indicates 1024 words have been written
                        next_state = S_FFT_IN_CONFIG;
                    else
                        next_state = S_DONE;
                end else
                    next_state = S_UART_WHO_AM_I_WAIT_BUSY_LOW;
            end
            
            
            // 9.
            
            S_FFT_IN_CONFIG: begin
                if (flit_transfer_counter_reg == 1024) //counter logic  // 1024 means 1024 (ALL) flits have been transferred
                    next_state = S_FFT_WAIT_TLAST;
                else
                    next_state = S_FFT_IN_ASSERT_TVALID;
            end
            
            S_FFT_IN_ASSERT_TVALID: begin  // both ready and valid need to be high for 1 clk cycle
                if (m_axis_data_tready) begin
                    next_state = S_FFT_IN_CONFIG; // input next flit
                end else
                    next_state = S_FFT_IN_ASSERT_TVALID; // stay in this state
            end
            
            
            // 10.
            
            /*S_FFT_WAIT_TVALID: begin
                if (s_axis_data_tvalid)
                    next_state = S_FIFO_OUT_WRITE_CONFIG;
                else
                    next_state = S_FFT_WAIT_TVALID;
            end
            
            S_FIFO_OUT_WRITE_CONFIG: begin
                next_state = S_FIFO_OUT_WRITE_ENABLE;
            end
            
            S_FIFO_OUT_WRITE_ENABLE: begin
                if (s_axis_data_tlast && s_axis_data_tvalid)
                    next_state = S_UART_FIFO_OUT_H_LATCH;
                else
                    next_state =  S_FIFO_OUT_WRITE_CONFIG;
            end*/
            
            S_FFT_WAIT_TLAST: begin
                // We can accept data if our buffer is not full
                s_axis_data_tready = !fifo_out_full;
                
                // We perform a write if the FFT has data AND we are ready
                if (s_axis_data_tvalid && s_axis_data_tready) begin
                    fifo_out_write_en = 1'b1;
                end
                
                // We transition away only when the LAST transfer is complete
                if (s_axis_data_tlast && s_axis_data_tvalid && s_axis_data_tready)
                    next_state = S_UART_FIFO_OUT_H_LATCH;
                else
                    next_state = S_FFT_WAIT_TLAST;
            end
            
            
            // 11. higher byte
            
            S_UART_FIFO_OUT_H_LATCH: begin
                // Just wait 1 clock cycle to latch the higher byte to uart_tx's data_to_transmit_reg
                next_state = S_UART_FIFO_OUT_H_PULSE_ENABLE;
            end
            
            S_UART_FIFO_OUT_H_PULSE_ENABLE: begin
                uart_tx_en_pulse_sig = !uart_busy_sig && rst_n;         // HIGH only when the UART TX module is NOT busy and NOT in reset
                // uart_tx_en_pulse_sig is HIGH for 1 cycle, since the FSM states last 1 clock cycle each
                
                if (uart_tx_en_pulse_sig)
                    next_state = S_UART_FIFO_OUT_H_WAIT_BUSY_LOW;     // Only transition to the next state once enable signal is HIGH
                else
                    next_state = S_UART_FIFO_OUT_H_PULSE_ENABLE;
            end
            
            S_UART_FIFO_OUT_H_WAIT_BUSY_LOW: begin
                // Transition when UART TX module is not busy, else wait here till communication is finished
                if (!uart_busy_sig)
                    next_state = S_UART_FIFO_OUT_L_LATCH;
                else
                    next_state = S_UART_FIFO_OUT_H_WAIT_BUSY_LOW;
            end
            
            
            // 12. lower byte
            
            S_UART_FIFO_OUT_L_LATCH: begin
                // Just wait 1 clock cycle to latch the lower byte to uart_tx's data_to_transmit_reg
                next_state = S_UART_FIFO_OUT_L_PULSE_ENABLE;
            end
            
            S_UART_FIFO_OUT_L_PULSE_ENABLE: begin
                uart_tx_en_pulse_sig = !uart_busy_sig && rst_n;         // HIGH only when the UART TX module is NOT busy and NOT in reset
                // uart_tx_en_pulse_sig is HIGH for 1 cycle, since the FSM states last 1 clock cycle each
                
                if (uart_tx_en_pulse_sig)
                    next_state = S_UART_FIFO_OUT_L_WAIT_BUSY_LOW;     // Only transition to the next state once enable signal is HIGH
                else
                    next_state = S_UART_FIFO_OUT_L_PULSE_ENABLE;
            end
            
            S_UART_FIFO_OUT_L_WAIT_BUSY_LOW: begin
                // Transition when UART TX module is not busy, else wait here till communication is finished
                if (!uart_busy_sig) begin
                    if (fifo_out_empty)
                        next_state = S_DONE;
                    else
                        next_state = S_UART_FIFO_OUT_H_LATCH;
                end else
                    next_state = S_UART_FIFO_OUT_L_WAIT_BUSY_LOW;
            end
            
            
            S_DONE: begin
                next_state = S_I2C_ACCEL_XOUT_CONFIG;    // Loop back to burst reading accelerometer values
            end
            
        endcase
    end
    
endmodule
